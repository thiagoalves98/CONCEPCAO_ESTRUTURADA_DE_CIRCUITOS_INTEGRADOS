library verilog;
use verilog.vl_types.all;
entity tristate_tb is
end tristate_tb;
