library verilog;
use verilog.vl_types.all;
entity mux8_tb is
end mux8_tb;
