library verilog;
use verilog.vl_types.all;
entity signextend_tb is
end signextend_tb;
