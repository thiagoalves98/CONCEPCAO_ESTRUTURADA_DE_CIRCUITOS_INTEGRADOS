library verilog;
use verilog.vl_types.all;
entity shiftleft2_tb is
end shiftleft2_tb;
