library verilog;
use verilog.vl_types.all;
entity flopr32_tb is
end flopr32_tb;
