library verilog;
use verilog.vl_types.all;
entity flopenr32_tb is
end flopenr32_tb;
