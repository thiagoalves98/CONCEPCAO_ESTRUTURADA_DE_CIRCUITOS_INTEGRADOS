module inversor_5(input logic a, output logic  y);
       
assign y = ~a;
	   
endmodule
