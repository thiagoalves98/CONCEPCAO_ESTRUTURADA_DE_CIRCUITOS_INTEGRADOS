library verilog;
use verilog.vl_types.all;
entity decoder5_32 is
    port(
        a               : in     vl_logic_vector(0 to 4);
        y_31_0          : out    vl_logic;
        y_30_0          : out    vl_logic;
        y_29_0          : out    vl_logic;
        y_28_0          : out    vl_logic;
        y_27_0          : out    vl_logic;
        y_26_0          : out    vl_logic;
        y_25_0          : out    vl_logic;
        y_24_0          : out    vl_logic;
        y_23_0          : out    vl_logic;
        y_22_0          : out    vl_logic;
        y_21_0          : out    vl_logic;
        y_20_0          : out    vl_logic;
        y_19_0          : out    vl_logic;
        y_18_0          : out    vl_logic;
        y_17_0          : out    vl_logic;
        y_16_0          : out    vl_logic;
        y_15_0          : out    vl_logic;
        y_14_0          : out    vl_logic;
        y_13_0          : out    vl_logic;
        y_12_0          : out    vl_logic;
        y_11_0          : out    vl_logic;
        y_10_0          : out    vl_logic;
        y_9_0           : out    vl_logic;
        y_8_0           : out    vl_logic;
        y_7_0           : out    vl_logic;
        y_6_0           : out    vl_logic;
        y_5_0           : out    vl_logic;
        y_4_0           : out    vl_logic;
        y_3_0           : out    vl_logic;
        y_2_0           : out    vl_logic;
        y_1_0           : out    vl_logic;
        y_0_0           : out    vl_logic
    );
end decoder5_32;
