library verilog;
use verilog.vl_types.all;
entity bank_tb is
end bank_tb;
