library verilog;
use verilog.vl_types.all;
entity controle_tb is
end controle_tb;
