library verilog;
use verilog.vl_types.all;
entity decoder5_32_tb is
end decoder5_32_tb;
