library verilog;
use verilog.vl_types.all;
entity shiftpc_tb is
end shiftpc_tb;
