library verilog;
use verilog.vl_types.all;
entity mux32_tb is
end mux32_tb;
