module mux32(input logic [0:4]s, input logic [0:31][0:0]d, output logic y); 

	logic y0, y1, y2, y3, y4, y5, y6, y7, y8, y9;

	//S -> 1 barramento de 4bits  [0:0][0:4]s ou implicitamente [0:4]s
	//D -> 32 barramentos de 1bit [0:31][0:0]d
	mux4 m1(d[0] [0:0], d[1] [0:0], d[2] [0:0], d[3] [0:0], s[0], s[1], y0);
	mux4 m2(d[4] [0:0], d[5] [0:0], d[6] [0:0], d[7] [0:0], s[0], s[1], y1);
	mux4 m3(d[8] [0:0], d[9] [0:0], d[10][0:0], d[11][0:0], s[0], s[1], y2);
	mux4 m4(d[12][0:0], d[13][0:0], d[14][0:0], d[15][0:0], s[0], s[1], y3);
	mux4 m5(d[16][0:0], d[17][0:0], d[18][0:0], d[19][0:0], s[0], s[1], y4);
	mux4 m6(d[20][0:0], d[21][0:0], d[22][0:0], d[23][0:0], s[0], s[1], y5);
	mux4 m7(d[24][0:0], d[25][0:0], d[26][0:0], d[27][0:0], s[0], s[1], y6);
	mux4 m8(d[28][0:0], d[29][0:0], d[30][0:0], d[31][0:0], s[0], s[1], y7);
	
	mux4 m9 (y0, y1, y2, y3, s[2], s[3], y8);
	mux4 m10(y4, y5, y6, y7, s[2], s[3], y9);
	
	mux2 m11(y8, y9, s[4], y);

endmodule
